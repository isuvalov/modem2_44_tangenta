library IEEE;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.std_logic_arith.all;


entity RScoder_ver2 is
	generic(R : natural := 16; --���-�� ����������� ����	   
			AmountByte: natural := 188 -- ���-�� ���� �� �����
			);	   
	 port(
		 reset: in std_logic;
		 clk : in STD_LOGIC;
		 CE : in STD_LOGIC;
		 StartOfCodePocket: out std_logic;
		 EndOfCodePocket: out std_logic;
		 PrevEndOfCodePocket: out std_logic;
		 EndAndStartOfCodePocket: out std_logic;		 
		 ByteIn : in STD_LOGIC_VECTOR(7 downto 0);
		 Ready : out STD_LOGIC;  --���������� ����� �������������� ����� ������ ???
		 CanGetData : out STD_LOGIC;	--���������� ����� ����� ���� ����������� ���� ������
		 ByteOut : out STD_LOGIC_VECTOR(7 downto 0)
	     );
end RScoder_ver2;


architecture RScoder_ver2 of RScoder_ver2 is

type TIntArray is array (0 to 238) of Integer;
type TG_matrix is array (1 to R) of TIntArray;
CONSTANT G_matrix:TG_matrix:=(
(169,44,125,233,138,206,215,201,16,197,254,6,125,194,58,12,126,147,218,99,33,187,205,44,60,77,225,233,183,219,204,221,1,9,19,18,138,229,237,221,252,204,255,154,71,107,199,91,218,131,158,229,122,107,207,247,100,74,170,213,162,118,250,92,172,178,188,57,75,137,145,24,44,198,54,175,171,162,132,146,154,138,187,85,208,98,144,232,85,249,46,28,18,121,97,2,203,148,239,67,194,86,26,150,37,74,6,94,60,179,18,202,161,129,215,203,161,88,186,97,110,191,30,33,212,239,42,120,202,162,21,157,116,83,112,110,185,36,47,213,246,180,187,232,76,97,141,50,114,94,66,185,209,104,35,242,44,183,12,65,196,114,162,99,194,221,13,145,25,185,162,238,16,209,192,3,227,90,79,162,42,118,131,169,213,228,251,189,78,176,211,162,73,99,62,135,154,230,175,197,168,181,240,237,13,218,202,223,143,220,138,165,32,225,46,35,100,166,29,70,105,19,22,152,237,107,204,39,93,136,197,250,27,51,10,41,114,33,59),
(1,179,252,26,150,127,82,131,94,109,148,100,214,161,213,19,145,104,29,194,107,193,3,215,161,72,239,134,32,2,88,227,230,255,211,242,109,196,110,194,250,127,166,23,93,154,96,190,213,91,135,208,148,167,165,96,78,177,6,64,92,250,203,34,138,178,243,230,215,121,233,195,2,28,248,173,216,34,130,169,122,229,106,157,104,243,57,204,206,165,149,144,253,46,23,23,32,124,105,196,159,169,114,219,114,240,208,168,211,25,82,11,14,86,29,245,15,149,131,212,107,98,119,22,240,41,111,45,97,67,226,92,179,200,145,122,248,102,115,197,65,114,84,231,167,34,191,95,134,220,78,212,191,65,22,91,232,229,158,81,7,112,251,186,191,237,207,109,248,143,48,100,121,22,123,141,215,161,88,198,34,114,247,130,67,160,98,129,132,38,192,90,58,81,152,83,111,153,125,210,255,23,187,123,255,131,195,147,119,155,163,162,150,130,141,80,154,1,35,225,237,179,30,136,19,48,232,94,196,84,245,120,229,242,128,199,157,122,13),
(22,224,232,141,166,121,37,158,83,206,239,186,63,101,190,137,95,152,99,208,114,183,57,226,230,151,81,158,6,38,247,112,238,131,56,25,78,64,129,70,90,15,240,202,83,248,16,168,181,12,3,170,168,49,69,66,142,91,176,70,41,120,76,32,13,51,77,251,254,124,106,81,34,133,95,192,161,177,216,134,197,198,57,228,228,168,237,69,66,111,94,25,90,146,249,13,193,10,35,25,119,6,11,66,95,103,222,33,153,103,211,137,117,205,12,203,139,208,68,84,72,131,244,199,91,175,230,13,246,8,170,173,98,19,194,13,188,113,144,51,47,214,174,40,220,112,189,200,79,119,161,136,160,13,235,200,186,104,185,244,204,23,25,54,9,151,188,220,216,62,230,98,180,13,191,108,142,18,141,49,9,6,171,225,194,99,27,144,160,39,72,169,88,247,122,117,63,85,161,237,201,101,211,254,42,244,88,241,22,82,39,233,31,143,121,39,190,199,128,106,94,42,77,104,205,182,197,118,184,98,196,67,215,159,128,88,215,45,104),
(176,77,2,71,4,141,147,11,80,167,170,130,88,206,157,100,211,23,192,69,57,220,36,98,119,75,95,254,234,54,221,170,24,225,245,38,144,59,82,220,242,161,3,183,208,18,220,30,240,51,246,118,77,233,114,46,97,38,83,138,41,20,161,71,69,172,152,13,59,207,228,195,10,110,167,130,160,206,50,248,193,76,104,61,11,170,88,42,65,35,228,74,7,5,100,41,243,140,200,132,232,203,127,150,22,247,10,5,180,80,121,69,94,35,39,242,28,61,22,178,192,91,71,29,149,153,153,209,155,153,19,232,64,11,67,86,115,128,146,170,48,227,120,105,237,42,252,34,72,148,184,223,15,89,52,85,147,206,178,206,104,76,120,63,199,84,37,36,29,166,81,76,172,51,44,7,116,232,111,226,7,52,128,27,219,223,210,216,133,209,112,39,185,126,178,65,50,242,136,85,53,109,11,193,76,114,98,213,173,35,219,77,104,215,4,64,4,108,187,242,251,40,137,218,122,140,77,65,21,225,150,29,82,32,40,14,216,62,189),
(250,193,226,132,89,168,2,43,20,167,42,3,45,187,9,210,17,238,106,88,198,187,170,85,12,249,76,217,51,42,253,180,23,36,36,141,56,89,115,59,54,57,145,2,223,201,130,228,99,210,252,63,205,84,248,195,162,251,6,187,43,221,87,141,206,251,58,133,42,255,149,122,178,39,230,244,31,1,248,178,249,223,206,120,166,46,77,99,58,216,53,180,50,102,250,3,246,218,163,110,103,34,50,49,219,140,94,65,107,183,40,27,62,27,172,248,137,254,2,233,216,140,108,196,72,186,65,69,179,58,245,6,123,249,86,41,179,131,43,122,166,39,97,67,90,18,32,186,24,3,143,93,249,204,189,246,36,94,129,115,132,82,237,224,220,174,166,127,7,248,7,195,83,138,183,246,103,241,1,206,58,243,22,122,243,175,33,249,140,92,144,209,103,33,119,94,64,33,161,127,18,159,200,67,51,49,16,108,184,121,61,110,115,111,193,224,204,107,129,110,140,62,158,239,146,99,71,103,208,108,22,213,89,169,198,42,52,91,68),
(139,133,30,185,171,171,48,49,31,48,9,175,220,200,117,30,193,84,37,30,116,241,133,213,30,143,184,23,249,188,80,247,240,73,220,152,162,116,15,121,29,76,211,138,19,177,101,176,47,18,196,176,33,163,226,8,118,224,188,22,230,34,126,164,79,167,13,56,131,201,50,187,5,90,254,232,247,66,177,249,169,214,232,99,33,150,167,82,206,85,47,22,8,224,154,114,184,114,4,191,139,6,132,62,16,153,9,37,10,70,11,215,138,199,131,23,105,119,141,254,206,226,39,64,144,150,64,215,186,238,71,47,135,83,117,113,150,214,48,59,206,74,16,126,132,166,252,244,190,99,91,48,64,91,104,4,137,4,73,21,19,128,15,153,5,214,253,107,21,184,165,157,247,78,231,123,63,17,250,92,52,51,130,157,106,251,72,147,182,109,201,205,95,19,226,11,69,192,47,133,176,186,174,158,16,248,206,146,10,246,86,161,6,50,152,101,85,156,12,212,136,116,143,13,185,252,25,238,208,119,72,181,55,201,59,240,46,24,209),
(212,17,33,180,60,51,181,165,160,47,6,213,11,225,31,208,212,194,62,10,240,142,7,31,222,20,227,18,72,66,155,55,38,231,182,242,29,173,189,104,240,58,171,199,249,250,62,34,218,189,101,203,25,200,234,195,42,113,90,29,106,234,119,52,194,162,80,180,238,104,117,101,33,91,40,246,131,139,221,99,237,44,44,181,112,223,251,220,15,245,112,27,56,207,112,37,88,182,4,20,130,184,238,53,179,23,69,252,46,54,104,240,197,167,217,169,5,64,92,29,165,87,105,201,48,230,208,86,44,198,205,94,156,6,131,46,52,202,34,145,203,255,176,107,165,20,46,237,155,75,162,30,242,199,10,251,158,214,161,230,244,124,252,32,164,98,162,65,237,80,196,2,12,53,204,137,168,169,164,134,26,56,161,86,60,180,127,110,247,228,16,181,164,112,167,19,31,36,200,31,128,80,150,103,234,122,3,22,165,188,115,39,158,106,23,201,71,74,121,174,130,119,57,36,196,80,219,43,117,234,71,29,140,247,176,19,159,192,30),
(178,187,78,64,195,224,252,51,88,174,233,66,138,95,55,151,173,176,155,40,243,131,112,104,141,155,133,130,233,15,162,152,41,200,56,119,133,244,180,190,146,16,226,33,78,31,200,194,123,67,79,140,206,255,10,194,143,53,225,169,125,231,84,209,224,95,139,164,181,187,48,120,10,13,5,222,120,227,72,167,233,154,95,100,32,120,153,132,148,147,166,5,218,31,229,76,159,102,147,245,64,232,137,236,180,172,83,223,110,173,247,204,178,96,104,99,235,219,45,118,157,174,30,144,36,21,205,233,242,76,93,29,239,144,207,3,97,171,135,209,167,18,140,207,48,143,57,8,24,1,164,237,149,54,2,68,148,101,94,108,246,1,28,234,116,167,244,250,82,162,48,255,255,135,93,238,36,74,208,196,173,151,161,19,165,203,20,72,9,86,83,112,136,178,222,70,153,212,210,198,179,71,34,143,241,179,222,60,7,184,203,73,192,15,57,210,133,95,33,238,116,93,206,143,61,34,176,102,147,62,228,249,50,180,59,185,230,102,8),
(33,207,116,85,100,253,22,250,179,62,13,217,141,212,146,87,64,65,46,164,61,66,165,13,149,223,192,158,83,127,33,4,144,97,80,168,83,254,207,18,13,188,187,70,35,49,105,42,92,23,199,52,123,177,201,225,197,229,12,7,208,234,100,142,216,25,214,94,198,137,71,240,5,116,160,20,239,1,183,172,3,205,43,205,170,23,140,138,22,15,254,70,149,53,48,245,90,75,77,177,171,202,56,77,217,222,156,153,34,159,61,233,173,206,150,126,2,17,98,2,33,12,94,11,126,15,88,42,247,139,228,193,154,77,55,152,162,92,206,97,50,110,163,159,149,31,147,180,191,210,43,5,43,242,51,193,57,69,5,108,2,65,120,35,180,210,207,8,50,243,219,19,127,57,201,69,165,206,8,169,137,58,251,128,245,214,64,149,2,224,128,42,2,183,95,146,226,250,197,180,239,114,148,25,231,111,173,104,48,169,156,138,84,155,98,60,213,220,183,43,129,236,237,122,180,66,12,149,180,167,88,103,33,183,228,110,14,243,163),
(72,63,63,147,60,20,189,40,24,74,117,224,41,58,197,85,95,25,101,160,222,204,202,187,241,94,73,39,168,212,84,75,167,66,123,233,193,115,175,165,2,38,84,48,167,220,147,173,14,231,42,231,138,132,98,80,33,64,85,23,198,169,23,238,211,251,166,63,120,87,139,212,238,4,162,5,7,46,244,77,39,106,60,115,195,135,182,200,210,19,74,219,255,211,224,107,144,77,65,26,6,11,2,116,129,92,51,77,101,162,38,251,208,77,142,243,71,62,67,183,232,102,114,36,179,116,252,189,236,54,124,33,227,47,217,221,50,205,186,213,91,252,159,231,247,64,56,243,123,110,38,129,168,44,211,191,223,15,130,9,54,205,128,246,148,222,182,205,56,152,50,114,241,210,213,49,136,194,94,201,90,240,129,179,155,118,136,92,166,122,22,65,87,140,16,82,25,58,95,60,95,130,165,197,125,195,169,156,20,249,192,19,83,194,222,67,252,162,90,245,143,155,227,61,43,75,105,155,188,134,94,165,12,226,157,239,161,116,65),
(188,171,116,14,36,31,32,68,76,202,197,238,171,33,38,238,221,255,71,227,41,132,44,41,60,22,93,120,86,183,117,208,10,212,229,157,94,219,91,43,168,163,232,135,103,19,140,139,243,202,45,48,118,62,230,158,12,28,63,227,90,124,63,213,10,250,123,121,67,12,117,221,55,255,51,133,59,74,48,21,158,144,48,141,157,4,228,198,121,135,114,5,61,173,215,98,16,234,231,15,18,116,223,250,228,188,199,115,202,13,68,28,117,150,121,245,125,156,37,71,91,171,171,251,211,25,12,239,135,161,10,117,25,201,14,53,5,227,237,12,104,233,166,239,65,243,45,22,80,59,97,254,46,223,39,119,92,174,36,78,154,149,128,6,254,16,180,148,218,224,213,217,22,94,88,22,176,209,167,19,177,224,52,61,5,192,161,73,120,13,87,91,191,209,137,205,129,192,29,141,193,172,164,141,175,35,249,175,115,209,78,87,219,80,163,213,31,168,172,76,195,40,100,178,21,159,234,123,24,137,84,200,48,99,82,38,76,40,41),
(12,4,2,234,48,44,193,247,238,106,33,51,71,82,197,215,60,53,249,231,131,221,247,148,59,118,221,195,125,121,237,172,249,118,5,29,163,49,225,130,146,242,97,124,202,146,103,154,141,177,250,66,70,131,31,113,225,153,107,179,193,221,51,246,84,130,209,228,197,6,182,138,101,106,234,201,219,25,215,241,129,160,100,133,140,20,151,83,115,77,109,41,253,48,95,133,231,39,130,14,246,220,217,186,62,113,74,92,97,107,245,232,69,101,72,252,172,16,65,215,63,11,162,203,94,187,87,40,67,165,134,65,160,90,184,118,147,232,32,97,178,22,29,17,140,179,18,156,53,203,251,199,214,160,237,61,207,89,95,159,65,185,183,32,255,39,200,14,66,124,194,148,115,62,245,35,143,143,201,133,93,54,162,56,177,67,166,163,120,162,119,117,181,31,145,111,89,149,58,59,168,150,228,158,85,169,143,114,28,131,239,179,30,16,186,145,170,153,218,200,235,18,116,162,136,224,197,124,155,116,175,27,76,168,100,103,5,44,229),
(140,53,209,113,165,51,71,67,1,164,110,69,230,140,249,13,48,27,115,197,243,46,236,206,91,233,126,174,166,222,173,42,73,103,178,36,82,24,241,38,81,70,19,216,2,141,15,39,220,92,187,65,22,1,101,133,204,178,39,215,118,93,106,242,44,103,174,72,82,184,246,59,179,29,9,2,146,30,73,21,72,206,13,59,111,85,1,1,12,246,163,83,8,155,219,136,208,65,48,79,197,155,134,168,29,109,21,92,147,183,74,69,31,67,14,29,11,222,88,170,198,33,226,182,146,73,230,212,152,134,5,190,10,155,162,169,12,209,227,156,30,229,187,139,38,103,125,194,179,35,227,129,200,163,99,33,4,170,145,69,48,110,124,139,235,56,10,56,102,56,185,48,98,124,34,199,252,42,138,12,216,193,231,46,132,239,17,111,67,156,122,178,20,137,7,243,214,208,125,112,82,26,141,36,179,19,25,159,107,62,204,171,66,22,254,121,44,220,66,65,88,47,128,26,98,207,52,181,88,3,62,24,164,121,4,11,72,17,98),
(222,242,226,170,213,49,156,224,45,4,130,63,146,208,205,91,124,175,116,172,123,135,28,146,222,62,165,5,120,171,142,241,72,28,175,24,128,139,246,173,196,1,2,217,78,234,76,85,72,45,3,98,165,254,247,22,105,154,202,76,152,48,238,3,219,13,32,73,124,80,227,175,69,16,254,134,24,221,220,180,223,236,186,49,167,210,108,24,61,25,76,111,249,74,128,31,235,124,107,51,121,95,6,238,131,75,60,184,76,208,29,75,172,42,236,109,244,247,200,67,181,39,41,92,191,184,102,198,213,215,31,252,60,103,140,189,25,69,9,136,141,110,145,162,140,61,240,11,17,30,66,83,127,134,217,231,95,210,8,86,34,227,33,163,189,183,248,81,3,214,119,241,94,156,142,132,79,196,139,197,35,158,48,57,69,63,62,52,172,166,166,53,66,203,93,99,57,169,95,120,204,64,90,99,228,220,18,129,204,85,154,176,119,14,172,132,149,246,114,182,109,144,16,142,244,138,159,219,190,56,6,141,231,176,138,141,216,246,50),
(137,149,144,119,123,208,140,7,231,243,8,46,93,210,48,136,111,21,101,48,144,145,212,87,222,181,38,48,170,128,202,218,195,247,77,204,201,80,214,162,197,165,63,212,91,135,80,140,159,38,51,211,158,108,201,68,204,156,69,19,30,33,244,176,112,142,121,150,142,251,93,105,228,205,181,219,107,74,45,135,98,14,6,91,18,209,237,203,249,175,54,14,12,83,106,228,224,28,69,33,115,206,177,149,26,118,231,6,244,43,179,208,79,166,151,19,105,98,47,232,112,151,1,21,183,134,95,254,11,135,42,87,33,113,114,191,51,223,88,208,9,116,132,54,251,172,114,157,122,43,102,204,66,224,222,144,172,240,151,38,186,83,177,101,227,233,192,245,233,141,132,124,246,79,184,216,248,189,203,217,34,154,240,185,224,167,201,120,9,157,211,244,150,6,227,251,181,191,140,129,195,7,109,7,20,46,17,34,170,170,132,86,190,111,33,244,94,15,134,194,27,60,59,162,211,61,235,15,183,11,230,194,81,184,89,59,252,228,36),
(26,208,103,127,245,156,84,151,125,81,154,208,220,23,41,157,22,142,24,8,224,184,26,141,116,162,103,201,181,131,47,59,254,218,225,127,78,139,47,39,131,106,232,199,221,11,121,142,129,4,78,113,221,206,175,185,213,76,234,137,88,189,216,214,30,65,90,238,50,96,82,26,48,62,155,119,137,32,45,232,127,224,38,61,35,91,92,38,240,108,190,225,60,110,118,34,183,253,43,220,107,36,193,228,213,154,174,141,37,225,25,196,247,156,34,196,52,219,110,10,12,200,8,209,253,128,7,25,137,64,73,46,188,194,10,150,223,87,234,148,132,224,92,79,110,222,210,180,174,16,150,6,144,126,120,26,201,41,93,70,180,137,24,220,47,18,96,105,150,137,198,151,6,170,77,212,66,2,137,128,88,129,1,234,117,134,122,57,104,112,137,152,24,251,109,232,3,155,125,58,191,14,139,18,142,25,89,168,20,127,40,51,162,108,126,185,101,133,252,171,218,13,158,139,221,131,146,227,9,125,189,31,233,179,205,180,8,44,59)
);



function gf_mul(a,b:std_logic_vector(7 downto 0)) return std_logic_vector is
variable answ:std_logic_vector(7 downto 0);
variable c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14:std_logic;	
begin
 -- (a7*x7+a6*x6+...+a0)*(b7*x7+b6*x6+...+b0)=c14*x14+c13*x13+...+c0
 -- c14*x14+c13*x13+...+c0 mod x8+x4+x3+x2+1 = answ	  
 -- �.�. ��� ���� ���� ������� ��� ����� ������������ ������ ��������� ���� �������� ������� �� ������� � �������� ��� � answ
 c0:=a(0) and b(0);
 c1:=(a(0) and b(1)) xor (a(1) and b(0));
 c2:=(a(0) and b(2)) xor (a(1) and b(1)) xor (a(2) and b(0));
 c3:=(a(0) and b(3)) xor (a(1) and b(2)) xor (a(2) and b(1)) xor (a(3) and b(0));
 c4:=(a(0) and b(4)) xor (a(1) and b(3)) xor (a(2) and b(2)) xor (a(3) and b(1)) xor (a(4) and b(0));
 c5:=(a(0) and b(5)) xor (a(1) and b(4)) xor (a(2) and b(3)) xor (a(3) and b(2)) xor (a(4) and b(1)) xor (a(5) and b(0));
 c6:=(a(0) and b(6)) xor (a(1) and b(5)) xor (a(2) and b(4)) xor (a(3) and b(3)) xor (a(4) and b(2)) xor (a(5) and b(1)) xor (a(6) and b(0));
 c7:=(a(0) and b(7)) xor (a(1) and b(6)) xor (a(2) and b(5)) xor (a(3) and b(4)) xor (a(4) and b(3)) xor (a(5) and b(2)) xor (a(6) and b(1)) xor (a(7) and b(0));
 c8:=(a(1) and b(7)) xor (a(2) and b(6)) xor (a(3) and b(5)) xor (a(4) and b(4)) xor (a(5) and b(3)) xor (a(6) and b(2)) xor (a(7) and b(1));
 c9:=(a(2) and b(7)) xor (a(3) and b(6)) xor (a(4) and b(5)) xor (a(5) and b(4)) xor (a(6) and b(3)) xor (a(7) and b(2));
c10:=(a(3) and b(7)) xor (a(4) and b(6)) xor (a(5) and b(5)) xor (a(6) and b(4)) xor (a(7) and b(3));
c11:=(a(4) and b(7)) xor (a(5) and b(6)) xor (a(6) and b(5)) xor (a(7) and b(4));
c12:=(a(5) and b(7)) xor (a(6) and b(6)) xor (a(7) and b(5));
c13:=(a(6) and b(7)) xor (a(7) and b(6));
c14:=(a(7) and b(7));
answ(7):=c7 xor c13 xor c12 xor c11;
answ(6):=c6 xor c12 xor c11 xor c10;
answ(5):=c5 xor c11 xor c10 xor c9;
answ(4):=c4 xor c14 xor c10 xor c9 xor c8;
answ(3):=c3 xor c11 xor c9 xor c8 xor c12;
answ(2):=c2 xor c10 xor c8 xor c13 xor c12;
answ(1):=c1 xor c9 xor c13 xor c14;
answ(0):=c0 xor c8 xor c14 xor c13 xor c12;
return answ;
end gf_mul;


component pincounter is
	 generic(NumberOfPins : natural := 8);		
	 port(
		 clk : in STD_LOGIC;
		 start : in STD_LOGIC;
		 en : in STD_LOGIC;
		 now : out STD_LOGIC;
		 data : out STD_LOGIC_VECTOR(NumberOfPins-1 downto 0)
	     );
end component;

attribute ramstyle : string;
attribute ramstyle of G_matrix : constant is "M9K";


type TScalar is array (1 to R) of std_logic_vector(7 downto 0);
type IScalar is array (1 to R) of Integer;

signal ccc,cnt_w1,cnt,cnt2,cntV:std_logic_vector(7 downto 0):=(others=>'0');
signal ccc2:std_logic_vector(7 downto 0):=x"00";
signal canGetd:std_logic:='1';
signal canGetd_w2,canGetd_w1:std_logic:='0';
signal Scalar,ScalarTRIG:TScalar:=(others=>x"00");
signal ByteIn_p1,ByteIn_w1,ByteIn_w2,ByteIn_w3:std_logic_vector(7 downto 0):=(others=>'0');

signal scI:IScalar:=(others=>0); 


signal DataInTest:std_logic_vector(7 downto 0):=(others=>'0');
signal Addsign,CE_w1,CE_w2,CE_w3:std_logic:='0';
--signal MUXcnt:std_logic_vector(R downto 0);

signal canGetd_p1:std_logic;
signal muxcnt:std_logic_vector(3 downto 0);
signal calccnt,test_cnt:std_logic_vector(7 downto 0):=(others=>'0');

begin



process (clk) is
begin		
	if rising_edge(clk) then 	
		if canGetd='1' and canGetd_w1='0' then
			--DataInTest<=CONV_STD_LOGIC_VECTOR(AmountByte-1,8);
			DataInTest<=CONV_STD_LOGIC_VECTOR(3,8);
		elsif (canGetd)='1' and CE='1' then	
			DataInTest<=DataInTest+1;
		end if;
	end if;
end process;


Ready<='1';
CanGetData<=canGetd_p1;

process (clk) is
begin		
	if rising_edge(clk) then 

            CE_w1<=CE;		
			CE_w2<=CE_w1;
			CE_w3<=CE_w2;

			ByteIn_w1<=ByteIn;
			ByteIn_w2<=ByteIn_w1;
			ByteIn_w3<=ByteIn_w2;
--		if reset='1' then
		if CE='1' and CE_w1='0' then
			cnt<=(others=>'0');
--			CE_w1<='0';
			EndOfCodePocket<='0';
			StartOfCodePocket<='0';
			canGetd_p1<='0';
			canGetd<='0';
		else
			if unsigned(cnt)<(AmountByte+R) then
				cnt<=cnt+1;
			else
				cnt<=(others=>'0');
			end if;

			if cnt=CONV_STD_LOGIC_VECTOR(AmountByte+R,8) then 
				canGetd_p1<='1';
	    	elsif cnt=CONV_STD_LOGIC_VECTOR(AmountByte,8) then
				canGetd_p1<='0';
			end if;
			
			canGetd<=canGetd_p1;	  

			if cnt=CONV_STD_LOGIC_VECTOR(0+1,8) then
				EndOfCodePocket<='1';
			else
				EndOfCodePocket<='0';
			end if;		

			if cnt=CONV_STD_LOGIC_VECTOR(1+1,8)  then
				StartOfCodePocket<='1';
			else 
				StartOfCodePocket<='0';
			end if;	  

		end if; --#reset


		if CE='1' then		
			if cnt=x"01" then 
				ByteIn_p1<=ByteIn;
			end if;
			
			if cnt=CONV_STD_LOGIC_VECTOR(AmountByte-2,8) then 
				Addsign<='1';
			else 
				Addsign<='0';
			end if;

			canGetd_w1<=canGetd;
			canGetd_w2<=canGetd_w1;
			cnt_w1<=cnt;
		end if;
		
		end if;
end process;

cnt2<=cnt-14;

process (clk) is
begin		
	if rising_edge(clk) then	
		if reset='1' then
			Scalar<=(others=>x"00");
			calccnt<=conv_std_logic_vector(239,calccnt'Length);
		else --# reset			
			if CE_w2='1' then
				if unsigned(cnt)<=188 then
					for k in 1 To R loop
						Scalar(k)<=Scalar(k) xor GF_Mul(ByteIn_w2,CONV_STD_LOGIC_VECTOR(G_matrix(k)(CONV_INTEGER(51+cnt-1)),8) );
					end loop;
				end if;
				if unsigned(calccnt)<255 then
					calccnt<=calccnt+1;
				end if;
			else
				if ce_w3='1' then
					ScalarTRIG<=Scalar;
				end if;
				Scalar<=(others=>x"00");
				calccnt<=conv_std_logic_vector(239,calccnt'Length);
			end if;
		end if; --# reset
	end if;
end process;

cntV<=cnt-1;

MuxDataForOut:process (clk) is
begin		
	if rising_edge(clk) then
		if ce_w3='1' then
			ByteOut<=ByteIn_w3;
			muxcnt<=(others=>'0');
			test_cnt<=test_cnt+1;
		else --# ce
			if unsigned(muxcnt)<R-1 then
				muxcnt<=muxcnt+1;
			end if; --# muxcnt
			for i in 0 to R-1 loop
				if muxcnt=i then
					ByteOut<=ScalarTRIG(i+1);
				end if; --# i
			end loop;
		end if; --# ce
	end if;
end process;


end RScoder_ver2;
